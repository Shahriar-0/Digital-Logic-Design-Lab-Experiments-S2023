module detector(input clk, Clk_EN, rst, serIn,
                output serOut, serOutValid, inc_cnt, )