module detector(input clk, Clk_EN, rst, serIn, Co
                output serOut, serOutValid, inc_cnt, rst_cnt)