module adder(input [17:0] a,b, output [17:0] s);

assign s = a+b;

endmodule
