module Exponential(); 
		   
endmodule

