module memoryRomImplementation();
    (* romstyle = "M9K")(* ram_inital_file = "sine.mif" *) reg [7:0] mem [3:0];