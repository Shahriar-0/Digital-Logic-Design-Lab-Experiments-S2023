module Controller();

	
endmodule

