module FreqSelector #(parameter N = 9)
                     (sel, clk, rst, co);
    
    input [4:0] sel;
    input clr, clk, rst;
    output co;

    
endmodule
