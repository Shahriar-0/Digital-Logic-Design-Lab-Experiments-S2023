module Datapath();
		 
endmodule

