module accelerator_wrappers(input clk , rst, start, input [1:0] U, input [5:0] V,output done, output out);