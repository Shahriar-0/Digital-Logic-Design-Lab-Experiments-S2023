module top_tb();
    reg start, rst, clk;
    reg [4:0] V;
    reg [1:0] U;
    wire done, wr_req;
    wire [20:0] wr_data;
    
    always #5 clk = ~clk;

    

endmodule